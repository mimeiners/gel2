* BODE-DIAGRAMM REIHENSCHWINGKREIS
C1 vo 0 1u
R1 N001 vi 10
V1 vi 0 AC 1
L1 N001 vo 100m

* ANALYSIS
.ac dec 50 10 1MEG

.end
